`timescale 1ns / 1ps

module conv2_weights_memory(
    input  wire               clk,
    input  wire               rst,
    input  wire               start,
    input  wire        [3:0]  output_filter,
    input  wire        [4:0]  input_filter,
    output wire signed [15:0] w0, w1,
    output wire done
);
    reg signed [15:0] weights0 [0:9][0:19];
    reg signed [15:0] weights1 [0:9][0:19];
    
    initial begin
        weights0[0][0] <=  -1086; weights0[0][1] <=    109; weights0[0][2] <=   -649; weights0[0][3] <=   -403; weights0[0][4] <=   -968; weights0[0][5] <=     34; weights0[0][6] <=  -1109; weights0[0][7] <=    851; weights0[0][8] <=    -72; weights0[0][9] <=   -174; weights0[0][10] <=    -38; weights0[0][11] <=      3; weights0[0][12] <=      7; weights0[0][13] <=   -810; weights0[0][14] <=    -12; weights0[0][15] <=    523; weights0[0][16] <=     54; weights0[0][17] <=    934; weights0[0][18] <=   -152; weights0[0][19] <=    -78; 
        weights0[1][0] <=   -357; weights0[1][1] <=    -47; weights0[1][2] <=   -152; weights0[1][3] <=   -273; weights0[1][4] <=      4; weights0[1][5] <=     22; weights0[1][6] <=   -439; weights0[1][7] <=   -123; weights0[1][8] <=    -26; weights0[1][9] <=   -549; weights0[1][10] <=     10; weights0[1][11] <=   -281; weights0[1][12] <=   -309; weights0[1][13] <=   -206; weights0[1][14] <=     42; weights0[1][15] <=     64; weights0[1][16] <=    -57; weights0[1][17] <=   -416; weights0[1][18] <=    238; weights0[1][19] <=     80; 
        weights0[2][0] <=   1360; weights0[2][1] <=   -447; weights0[2][2] <=    -39; weights0[2][3] <=   -404; weights0[2][4] <=  -1291; weights0[2][5] <=    152; weights0[2][6] <=   1519; weights0[2][7] <=   -151; weights0[2][8] <=    488; weights0[2][9] <=   -858; weights0[2][10] <=   -190; weights0[2][11] <=    116; weights0[2][12] <=    103; weights0[2][13] <=   -575; weights0[2][14] <=    -91; weights0[2][15] <=     88; weights0[2][16] <=   -447; weights0[2][17] <=   -400; weights0[2][18] <=   1262; weights0[2][19] <=  -2028; 
        weights0[3][0] <=    -14; weights0[3][1] <=   -115; weights0[3][2] <=   -318; weights0[3][3] <=    -55; weights0[3][4] <=   -246; weights0[3][5] <=    -94; weights0[3][6] <=   -165; weights0[3][7] <=   -223; weights0[3][8] <=   -256; weights0[3][9] <=   -383; weights0[3][10] <=   -341; weights0[3][11] <=   -304; weights0[3][12] <=    205; weights0[3][13] <=   -222; weights0[3][14] <=   -298; weights0[3][15] <=    -63; weights0[3][16] <=     75; weights0[3][17] <=     17; weights0[3][18] <=   -195; weights0[3][19] <=   -283; 
        weights0[4][0] <=    403; weights0[4][1] <=    610; weights0[4][2] <=     24; weights0[4][3] <=    397; weights0[4][4] <=   -925; weights0[4][5] <=    -14; weights0[4][6] <=    299; weights0[4][7] <=  -1642; weights0[4][8] <=  -1716; weights0[4][9] <=    -42; weights0[4][10] <=     83; weights0[4][11] <=   -842; weights0[4][12] <=   -116; weights0[4][13] <=   1700; weights0[4][14] <=    147; weights0[4][15] <=  -1061; weights0[4][16] <=    -50; weights0[4][17] <=  -3414; weights0[4][18] <=    361; weights0[4][19] <=   -490; 
        weights0[5][0] <=   -469; weights0[5][1] <=    237; weights0[5][2] <=    -21; weights0[5][3] <=    513; weights0[5][4] <=   -388; weights0[5][5] <=     25; weights0[5][6] <=   -544; weights0[5][7] <=   -389; weights0[5][8] <=    113; weights0[5][9] <=    -21; weights0[5][10] <=   -331; weights0[5][11] <=    160; weights0[5][12] <=     94; weights0[5][13] <=   -339; weights0[5][14] <=   -135; weights0[5][15] <=    126; weights0[5][16] <=     81; weights0[5][17] <=   -114; weights0[5][18] <=    685; weights0[5][19] <=   -153; 
        weights0[6][0] <=   -336; weights0[6][1] <=    -42; weights0[6][2] <=   -231; weights0[6][3] <=   -263; weights0[6][4] <=    136; weights0[6][5] <=   -168; weights0[6][6] <=   -411; weights0[6][7] <=   -191; weights0[6][8] <=    -42; weights0[6][9] <=   -609; weights0[6][10] <=    123; weights0[6][11] <=   -630; weights0[6][12] <=   -499; weights0[6][13] <=   -807; weights0[6][14] <=    -43; weights0[6][15] <=   -255; weights0[6][16] <=   -622; weights0[6][17] <=   -565; weights0[6][18] <=     63; weights0[6][19] <=    113; 
        weights0[7][0] <=   -646; weights0[7][1] <=   -200; weights0[7][2] <=   1134; weights0[7][3] <=   -443; weights0[7][4] <=  -1376; weights0[7][5] <=   -239; weights0[7][6] <=   -755; weights0[7][7] <=   -930; weights0[7][8] <=   -145; weights0[7][9] <=   1344; weights0[7][10] <=     84; weights0[7][11] <=     46; weights0[7][12] <=   -171; weights0[7][13] <=  -3614; weights0[7][14] <=   -189; weights0[7][15] <=     79; weights0[7][16] <=    -24; weights0[7][17] <=   -877; weights0[7][18] <=   1105; weights0[7][19] <=   -118; 
        weights0[8][0] <=    578; weights0[8][1] <=    569; weights0[8][2] <=    833; weights0[8][3] <=    188; weights0[8][4] <=  -1058; weights0[8][5] <=    128; weights0[8][6] <=    942; weights0[8][7] <=  -2253; weights0[8][8] <=   -968; weights0[8][9] <=    741; weights0[8][10] <=   -395; weights0[8][11] <=   -321; weights0[8][12] <=   -160; weights0[8][13] <=    513; weights0[8][14] <=   -520; weights0[8][15] <=   -764; weights0[8][16] <=   -124; weights0[8][17] <=  -2933; weights0[8][18] <=    636; weights0[8][19] <=  -1162; 
        weights0[9][0] <=  -2197; weights0[9][1] <=   -417; weights0[9][2] <=    355; weights0[9][3] <=   -178; weights0[9][4] <=   -399; weights0[9][5] <=    -23; weights0[9][6] <=  -1846; weights0[9][7] <=     80; weights0[9][8] <=   -118; weights0[9][9] <=    262; weights0[9][10] <=   -118; weights0[9][11] <=    118; weights0[9][12] <=    245; weights0[9][13] <=   -573; weights0[9][14] <=      0; weights0[9][15] <=     69; weights0[9][16] <=   -193; weights0[9][17] <=   -194; weights0[9][18] <=   -519; weights0[9][19] <=    647; 
        
        weights1[0][0] <=    540; weights1[0][1] <=   -702; weights1[0][2] <=  -1561; weights1[0][3] <=   -292; weights1[0][4] <=   1121; weights1[0][5] <=   -113; weights1[0][6] <=    496; weights1[0][7] <=    762; weights1[0][8] <=    675; weights1[0][9] <=  -1965; weights1[0][10] <=     27; weights1[0][11] <=    843; weights1[0][12] <=   -103; weights1[0][13] <=    585; weights1[0][14] <=     34; weights1[0][15] <=   1161; weights1[0][16] <=    242; weights1[0][17] <=    408; weights1[0][18] <=   -257; weights1[0][19] <=     76; 
        weights1[1][0] <=   -251; weights1[1][1] <=    239; weights1[1][2] <=   -214; weights1[1][3] <=   -290; weights1[1][4] <=   -523; weights1[1][5] <=    421; weights1[1][6] <=   -187; weights1[1][7] <=   -146; weights1[1][8] <=   -600; weights1[1][9] <=   -257; weights1[1][10] <=     -9; weights1[1][11] <=   -602; weights1[1][12] <=   -499; weights1[1][13] <=   -115; weights1[1][14] <=     20; weights1[1][15] <=   -740; weights1[1][16] <=   -513; weights1[1][17] <=   -518; weights1[1][18] <=   -360; weights1[1][19] <=   -733; 
        weights1[2][0] <=    328; weights1[2][1] <=    -72; weights1[2][2] <=  -1184; weights1[2][3] <=   -112; weights1[2][4] <=    -59; weights1[2][5] <=    185; weights1[2][6] <=    444; weights1[2][7] <=    -26; weights1[2][8] <=   -461; weights1[2][9] <=  -1230; weights1[2][10] <=      6; weights1[2][11] <=   -361; weights1[2][12] <=   -146; weights1[2][13] <=   -388; weights1[2][14] <=    -13; weights1[2][15] <=   -411; weights1[2][16] <=   -245; weights1[2][17] <=    187; weights1[2][18] <=  -1319; weights1[2][19] <=   -588; 
        weights1[3][0] <=    -33; weights1[3][1] <=   -202; weights1[3][2] <=    -94; weights1[3][3] <=   -149; weights1[3][4] <=     13; weights1[3][5] <=    277; weights1[3][6] <=   -208; weights1[3][7] <=   -177; weights1[3][8] <=   -125; weights1[3][9] <=     54; weights1[3][10] <=    -52; weights1[3][11] <=    243; weights1[3][12] <=   -164; weights1[3][13] <=   -217; weights1[3][14] <=      2; weights1[3][15] <=   -268; weights1[3][16] <=   -207; weights1[3][17] <=     29; weights1[3][18] <=      8; weights1[3][19] <=     38; 
        weights1[4][0] <=     55; weights1[4][1] <=    -57; weights1[4][2] <=  -1580; weights1[4][3] <=    329; weights1[4][4] <=  -1889; weights1[4][5] <=    -56; weights1[4][6] <=    317; weights1[4][7] <=    325; weights1[4][8] <=    -97; weights1[4][9] <=   -633; weights1[4][10] <=   -238; weights1[4][11] <=    -64; weights1[4][12] <=     56; weights1[4][13] <=   -299; weights1[4][14] <=   -349; weights1[4][15] <=   -254; weights1[4][16] <=     -2; weights1[4][17] <=    149; weights1[4][18] <=   -105; weights1[4][19] <=  -2373; 
        weights1[5][0] <=     89; weights1[5][1] <=    508; weights1[5][2] <=    -38; weights1[5][3] <=    242; weights1[5][4] <=  -1651; weights1[5][5] <=   -104; weights1[5][6] <=     94; weights1[5][7] <=   1226; weights1[5][8] <=   -206; weights1[5][9] <=     38; weights1[5][10] <=    -72; weights1[5][11] <=  -3206; weights1[5][12] <=     61; weights1[5][13] <=  -1870; weights1[5][14] <=   -208; weights1[5][15] <=  -2848; weights1[5][16] <=     40; weights1[5][17] <=    998; weights1[5][18] <=    -69; weights1[5][19] <=  -3002; 
        weights1[6][0] <=   -204; weights1[6][1] <=     98; weights1[6][2] <=   -471; weights1[6][3] <=   -105; weights1[6][4] <=   -164; weights1[6][5] <=   -285; weights1[6][6] <=   -294; weights1[6][7] <=   -414; weights1[6][8] <=   -793; weights1[6][9] <=   -223; weights1[6][10] <=   -412; weights1[6][11] <=   -825; weights1[6][12] <=   -538; weights1[6][13] <=   -204; weights1[6][14] <=    -86; weights1[6][15] <=   -768; weights1[6][16] <=   -676; weights1[6][17] <=   -188; weights1[6][18] <=   -681; weights1[6][19] <=    -42; 
        weights1[7][0] <=  -1156; weights1[7][1] <=   -396; weights1[7][2] <=   -269; weights1[7][3] <=   -196; weights1[7][4] <=   -311; weights1[7][5] <=    226; weights1[7][6] <=   -406; weights1[7][7] <=    432; weights1[7][8] <=    354; weights1[7][9] <=   -822; weights1[7][10] <=     30; weights1[7][11] <=    511; weights1[7][12] <=   -309; weights1[7][13] <=   -263; weights1[7][14] <=   -403; weights1[7][15] <=    448; weights1[7][16] <=   -560; weights1[7][17] <=    501; weights1[7][18] <=  -2215; weights1[7][19] <=    280; 
        weights1[8][0] <=   -665; weights1[8][1] <=    247; weights1[8][2] <=  -2187; weights1[8][3] <=    -96; weights1[8][4] <=   -334; weights1[8][5] <=    318; weights1[8][6] <=  -1045; weights1[8][7] <=    605; weights1[8][8] <=    195; weights1[8][9] <=  -1376; weights1[8][10] <=    127; weights1[8][11] <=    317; weights1[8][12] <=   -196; weights1[8][13] <=   -458; weights1[8][14] <=    181; weights1[8][15] <=    139; weights1[8][16] <=    120; weights1[8][17] <=    -26; weights1[8][18] <=   -449; weights1[8][19] <=    -41; 
        weights1[9][0] <=    821; weights1[9][1] <=    -47; weights1[9][2] <=  -1626; weights1[9][3] <=   -120; weights1[9][4] <=    109; weights1[9][5] <=     -0; weights1[9][6] <=   1056; weights1[9][7] <=    243; weights1[9][8] <=    626; weights1[9][9] <=  -1808; weights1[9][10] <=   -234; weights1[9][11] <=    256; weights1[9][12] <=   -170; weights1[9][13] <=   -201; weights1[9][14] <=    237; weights1[9][15] <=    714; weights1[9][16] <=   -272; weights1[9][17] <=    125; weights1[9][18] <=   -305; weights1[9][19] <=    -67;
    end
    
    assign w0   = weights0[output_filter][input_filter];
    assign w1   = weights1[output_filter][input_filter];
    assign done = (start == 1) ? 1 : 0;
endmodule
