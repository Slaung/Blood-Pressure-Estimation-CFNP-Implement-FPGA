`timescale 1ns / 1ps

module fr_weights_memory(
    input  wire                clk,
    input  wire                rst,
    input  wire                start,
    input  wire        [ 2: 0] output_filter_m,
    input  wire        [ 2: 0] output_filter_v,
    input  wire        [ 4: 0] input_filter,
    output wire signed [15: 0] m,
    output wire signed [15: 0] v,
    output wire                done
);
    reg signed [15:0] wm [0:4][0:20];
    reg signed [15:0] wv [0:4][0:20];

    initial begin
        wm[0][0] <=   463; wm[0][1] <=  -312; wm[0][2] <=  -243; wm[0][3] <=    46; wm[0][4] <=   374; wm[0][5] <=  -339; wm[0][6] <=    75; wm[0][7] <=   401; wm[0][8] <=  -120; wm[0][9] <=   356; wm[0][10] <=    61; wm[0][11] <=  -338; wm[0][12] <=   513; wm[0][13] <=   324; wm[0][14] <=   -84; wm[0][15] <=   382; wm[0][16] <=   224; wm[0][17] <=   -95; wm[0][18] <=  -282; wm[0][19] <=   410; wm[0][20] <=    97; 
        wm[1][0] <=   458; wm[1][1] <=  -309; wm[1][2] <=  -249; wm[1][3] <=    48; wm[1][4] <=   376; wm[1][5] <=  -323; wm[1][6] <=    76; wm[1][7] <=   409; wm[1][8] <=  -113; wm[1][9] <=   352; wm[1][10] <=    83; wm[1][11] <=  -327; wm[1][12] <=   505; wm[1][13] <=   343; wm[1][14] <=   -78; wm[1][15] <=   378; wm[1][16] <=   243; wm[1][17] <=   -81; wm[1][18] <=  -271; wm[1][19] <=   413; wm[1][20] <=   108; 
        wm[2][0] <=   459; wm[2][1] <=  -311; wm[2][2] <=  -244; wm[2][3] <=    42; wm[2][4] <=   370; wm[2][5] <=  -339; wm[2][6] <=    73; wm[2][7] <=   402; wm[2][8] <=  -120; wm[2][9] <=   355; wm[2][10] <=    62; wm[2][11] <=  -338; wm[2][12] <=   511; wm[2][13] <=   324; wm[2][14] <=   -84; wm[2][15] <=   381; wm[2][16] <=   225; wm[2][17] <=   -94; wm[2][18] <=  -283; wm[2][19] <=   410; wm[2][20] <=    98; 
        wm[3][0] <=   457; wm[3][1] <=  -309; wm[3][2] <=  -249; wm[3][3] <=    48; wm[3][4] <=   376; wm[3][5] <=  -323; wm[3][6] <=    76; wm[3][7] <=   410; wm[3][8] <=  -114; wm[3][9] <=   352; wm[3][10] <=    83; wm[3][11] <=  -328; wm[3][12] <=   505; wm[3][13] <=   342; wm[3][14] <=   -79; wm[3][15] <=   378; wm[3][16] <=   242; wm[3][17] <=   -82; wm[3][18] <=  -271; wm[3][19] <=   412; wm[3][20] <=   107; 
        wm[4][0] <=   463; wm[4][1] <=  -311; wm[4][2] <=  -242; wm[4][3] <=    46; wm[4][4] <=   374; wm[4][5] <=  -339; wm[4][6] <=    76; wm[4][7] <=   401; wm[4][8] <=  -120; wm[4][9] <=   356; wm[4][10] <=    60; wm[4][11] <=  -339; wm[4][12] <=   513; wm[4][13] <=   324; wm[4][14] <=   -85; wm[4][15] <=   382; wm[4][16] <=   224; wm[4][17] <=   -95; wm[4][18] <=  -282; wm[4][19] <=   410; wm[4][20] <=    97; 
        
        wv[0][0] <=    23; wv[0][1] <=    69; wv[0][2] <=    84; wv[0][3] <=    38; wv[0][4] <=    25; wv[0][5] <=     6; wv[0][6] <=    58; wv[0][7] <=     4; wv[0][8] <=    43; wv[0][9] <=    30; wv[0][10] <=     1; wv[0][11] <=    14; wv[0][12] <=    14; wv[0][13] <=     2; wv[0][14] <=    56; wv[0][15] <=     6; wv[0][16] <=     3; wv[0][17] <=     4; wv[0][18] <=     2; wv[0][19] <=     2; wv[0][20] <=    77; 
        wv[1][0] <=    25; wv[1][1] <=    88; wv[1][2] <=   129; wv[1][3] <=    56; wv[1][4] <=    34; wv[1][5] <=     7; wv[1][6] <=    91; wv[1][7] <=     5; wv[1][8] <=    51; wv[1][9] <=    38; wv[1][10] <=     2; wv[1][11] <=    15; wv[1][12] <=    16; wv[1][13] <=     2; wv[1][14] <=    72; wv[1][15] <=     7; wv[1][16] <=     3; wv[1][17] <=     5; wv[1][18] <=     3; wv[1][19] <=     3; wv[1][20] <=    95; 
        wv[2][0] <=    24; wv[2][1] <=    69; wv[2][2] <=    78; wv[2][3] <=    48; wv[2][4] <=    31; wv[2][5] <=     6; wv[2][6] <=    59; wv[2][7] <=     4; wv[2][8] <=    48; wv[2][9] <=    31; wv[2][10] <=     2; wv[2][11] <=    14; wv[2][12] <=    14; wv[2][13] <=     2; wv[2][14] <=    69; wv[2][15] <=     6; wv[2][16] <=     3; wv[2][17] <=     4; wv[2][18] <=     2; wv[2][19] <=     3; wv[2][20] <=    73; 
        wv[3][0] <=    25; wv[3][1] <=    84; wv[3][2] <=   128; wv[3][3] <=    57; wv[3][4] <=    35; wv[3][5] <=     7; wv[3][6] <=    92; wv[3][7] <=     5; wv[3][8] <=    52; wv[3][9] <=    39; wv[3][10] <=     2; wv[3][11] <=    15; wv[3][12] <=    16; wv[3][13] <=     2; wv[3][14] <=    74; wv[3][15] <=     7; wv[3][16] <=     3; wv[3][17] <=     5; wv[3][18] <=     3; wv[3][19] <=     3; wv[3][20] <=   101; 
        wv[4][0] <=    23; wv[4][1] <=    68; wv[4][2] <=    86; wv[4][3] <=    38; wv[4][4] <=    25; wv[4][5] <=     6; wv[4][6] <=    56; wv[4][7] <=     4; wv[4][8] <=    44; wv[4][9] <=    30; wv[4][10] <=     1; wv[4][11] <=    14; wv[4][12] <=    14; wv[4][13] <=     2; wv[4][14] <=    57; wv[4][15] <=     6; wv[4][16] <=     2; wv[4][17] <=     4; wv[4][18] <=     2; wv[4][19] <=     3; wv[4][20] <=    76; 
    end

    assign m    = (start == 1)? wm[output_filter_m][input_filter] : 0;
    assign v    = (start == 1)? wv[output_filter_v][input_filter] : 0;
    assign done = (start == 1)? 1 : 0;
endmodule